magic
tech scmos
timestamp 1638744199
<< nwell >>
rect 2 0 26 20
rect 32 0 88 20
rect 2 -50 26 -30
<< ntransistor >>
rect 13 -12 15 -8
rect 13 -62 15 -58
rect 44 -62 46 -58
rect 54 -62 56 -58
rect 64 -62 66 -58
rect 74 -62 76 -58
<< ptransistor >>
rect 13 6 15 14
rect 44 6 46 14
rect 54 6 56 14
rect 64 6 66 14
rect 74 6 76 14
rect 13 -44 15 -36
<< ndiffusion >>
rect 12 -12 13 -8
rect 15 -12 16 -8
rect 12 -62 13 -58
rect 15 -62 16 -58
rect 42 -62 44 -58
rect 46 -62 54 -58
rect 56 -62 58 -58
rect 62 -62 64 -58
rect 66 -62 74 -58
rect 76 -62 78 -58
<< pdiffusion >>
rect 12 6 13 14
rect 15 6 16 14
rect 42 6 44 14
rect 46 6 54 14
rect 56 6 58 14
rect 62 6 64 14
rect 66 6 74 14
rect 76 6 78 14
rect 12 -44 13 -36
rect 15 -44 16 -36
<< ndcontact >>
rect 8 -12 12 -8
rect 16 -12 20 -8
rect 8 -62 12 -58
rect 16 -62 20 -58
rect 38 -62 42 -58
rect 58 -62 62 -58
rect 78 -62 82 -58
<< pdcontact >>
rect 8 6 12 14
rect 16 6 20 14
rect 38 6 42 14
rect 58 6 62 14
rect 78 6 82 14
rect 8 -44 12 -36
rect 16 -44 20 -36
<< polysilicon >>
rect 44 24 86 26
rect 13 14 15 17
rect 44 14 46 24
rect 54 14 56 17
rect 64 14 66 17
rect 74 14 76 17
rect 13 -8 15 6
rect 44 -5 46 6
rect 54 -9 56 6
rect 44 -11 56 -9
rect 13 -15 15 -12
rect 13 -36 15 -33
rect 13 -58 15 -44
rect 44 -58 46 -11
rect 64 -14 66 6
rect 54 -16 66 -14
rect 54 -58 56 -16
rect 74 -48 76 6
rect 64 -50 76 -48
rect 64 -58 66 -50
rect 84 -53 86 24
rect 74 -55 86 -53
rect 74 -58 76 -55
rect 13 -65 15 -62
rect 44 -78 46 -62
rect 54 -65 56 -62
rect 64 -86 66 -62
rect 74 -65 76 -62
<< polycontact >>
rect 9 -5 13 -1
rect 40 -5 44 -1
rect 9 -55 13 -51
rect 50 -25 54 -21
rect 40 -78 44 -74
rect 60 -86 64 -82
<< metal1 >>
rect -21 20 88 24
rect -21 -5 -17 -1
rect -7 -26 -3 20
rect 8 14 12 20
rect 38 14 42 20
rect 78 14 82 20
rect 16 -1 20 6
rect 5 -5 9 -1
rect 16 -5 40 -1
rect 16 -8 20 -5
rect 8 -16 12 -12
rect 2 -20 35 -16
rect -7 -30 26 -26
rect 8 -36 12 -30
rect 16 -51 20 -44
rect -21 -55 -8 -51
rect -3 -55 9 -51
rect 16 -55 23 -51
rect 16 -58 20 -55
rect 8 -66 12 -62
rect 31 -66 35 -20
rect 43 -25 50 -21
rect 58 -27 62 6
rect 58 -31 90 -27
rect 58 -58 62 -31
rect 38 -66 42 -62
rect 78 -66 82 -62
rect -21 -70 88 -66
rect -2 -78 40 -74
rect 29 -86 60 -82
<< m2contact >>
rect -17 -6 -12 -1
rect 0 -6 5 -1
rect -8 -56 -3 -51
rect 23 -56 28 -51
rect 38 -26 43 -21
rect -7 -78 -2 -73
rect 24 -86 29 -81
<< metal2 >>
rect -12 -6 0 -2
rect -16 -21 -12 -6
rect -16 -25 38 -21
rect -7 -73 -3 -56
rect 24 -81 28 -56
<< labels >>
rlabel metal1 86 -31 90 -27 7 out
rlabel metal1 -21 -5 -17 -1 3 in1
rlabel metal1 -21 -55 -17 -51 3 in2
rlabel metal1 -21 -70 88 -66 1 gnd
rlabel metal1 -21 20 88 24 5 vdd
<< end >>